module MiniProject;
endmodule